library verilog;
use verilog.vl_types.all;
entity praca4_vlg_vec_tst is
end praca4_vlg_vec_tst;
