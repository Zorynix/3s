library verilog;
use verilog.vl_types.all;
entity praca5_vlg_vec_tst is
end praca5_vlg_vec_tst;
