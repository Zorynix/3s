library verilog;
use verilog.vl_types.all;
entity praca2kostya_vlg_vec_tst is
end praca2kostya_vlg_vec_tst;
