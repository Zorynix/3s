library verilog;
use verilog.vl_types.all;
entity praca5_vlg_check_tst is
    port(
        A_more_B        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end praca5_vlg_check_tst;
