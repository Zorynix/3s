library verilog;
use verilog.vl_types.all;
entity praca2tima_vlg_vec_tst is
end praca2tima_vlg_vec_tst;
