library verilog;
use verilog.vl_types.all;
entity practica1_vlg_vec_tst is
end practica1_vlg_vec_tst;
