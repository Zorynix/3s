library verilog;
use verilog.vl_types.all;
entity pract3_vlg_vec_tst is
end pract3_vlg_vec_tst;
