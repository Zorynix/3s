library verilog;
use verilog.vl_types.all;
entity praca4 is
    port(
        x0              : in     vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        Y0              : out    vl_logic;
        Y1              : out    vl_logic
    );
end praca4;
