library verilog;
use verilog.vl_types.all;
entity pr1timfad_vlg_vec_tst is
end pr1timfad_vlg_vec_tst;
