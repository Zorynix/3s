library verilog;
use verilog.vl_types.all;
entity praca6_vlg_vec_tst is
end praca6_vlg_vec_tst;
