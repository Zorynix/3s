library verilog;
use verilog.vl_types.all;
entity pract3 is
    port(
        Y0              : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic;
        Y1              : out    vl_logic
    );
end pract3;
