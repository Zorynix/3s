library verilog;
use verilog.vl_types.all;
entity praca5 is
    port(
        A_more_B        : out    vl_logic;
        A2              : in     vl_logic;
        B2              : in     vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        A0              : in     vl_logic;
        B0              : in     vl_logic
    );
end praca5;
