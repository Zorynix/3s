library verilog;
use verilog.vl_types.all;
entity pract2_vlg_vec_tst is
end pract2_vlg_vec_tst;
