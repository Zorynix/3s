library verilog;
use verilog.vl_types.all;
entity pract7_vlg_vec_tst is
end pract7_vlg_vec_tst;
